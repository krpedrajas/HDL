library ieee;
use ieee.std_logic_1164.all;

entity tb_tl is
end tb_tl;

architecture traffic_light of tb_tl is
    component tl is
    port(
        x : in std_logic_vector(2 downto 0);
        gyr : out std_logic_vector(5 downto 0)
    );
end component;

    signal tb_x : std_logic_vector(2 downto 0);
    signal tb_gyr : std_logic_vector(5 downto 0);

begin
    tl_module : tl port map(tb_x, tb_gyr);
    process
    begin
        tb_x <= "000";
        wait for 10 ns;

        tb_x <= "001";
        wait for 10 ns;

        tb_x <= "010";
        wait for 10 ns;

        tb_x <= "011";
        wait for 10 ns;

        tb_x <= "100";
        wait for 10 ns;

        tb_x <= "101";
        wait for 10 ns;

        wait;
    end process;
end traffic_light;